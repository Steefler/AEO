----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:41:45 10/21/2016 
-- Design Name: 
-- Module Name:    top - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity transform is
    Port ( switches : in  STD_LOGIC_VECTOR (7 downto 0);
           data : out  STD_LOGIC_VECTOR (15 downto 0));
end transform;

architecture Behavioral of transform is

begin

PROCESS(switches)
BEGIN
data <= "0000000000000000";

   IF (switches(6) = '1') THEN data (15 downto 12) <= "1111";
	END IF;
   IF (switches(4) = '1') THEN data (11 downto 8) <= "1111";
	END IF;
   IF (switches(2) = '1') THEN data (7 downto 4) <= "1111";
	END IF;
   IF (switches(0) = '1') THEN data (3 downto 0) <= "1111";
	END IF;

END PROCESS;


end Behavioral;

